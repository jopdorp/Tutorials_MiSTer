function int multiply(int a,b);
	return (a >>> 10) * (b >>> 10);
endfunction