function int divide(longint a, b);
	return (a <<< 10 )/ (b >>> 10);
endfunction