function int multiply(longint a,b);
	return (a * b) >>> 20;
endfunction