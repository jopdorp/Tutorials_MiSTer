function int divide(longint a, b);
	return (a <<< 20 )/ b;
endfunction